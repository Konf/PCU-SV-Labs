module my_module_name(

);

endmodule
