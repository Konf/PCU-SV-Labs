module xor_gate(
  input  logic a,
  input  logic b,
  output logic result
);

  assign result = a ^ b;

endmodule
