module stopwatch (
  input  logic clk,
  input  logic reset,
  input  logic start_stop,

  output logic [6:0] hex0,
  output logic [6:0] hex1,
  output logic [6:0] hex2,
  output logic [6:0] hex3
);

endmodule
