module not_gate(
  input  logic a,
  output logic result
);

  assign result = ~a;

endmodule
